module mul_param#(parameter n=32,m=8)(input [(n-1):0]a,b,
output reg [(n-1):0]out,
output reg overflow,underflow);
wire sign;
wire[m:0]expo_add;
wire[m+1:0]expo,temp;
wire[2*(n-m)-1:0] mant_mul;
wire[n-m-2:0]mant;
wire [(n-1):0]temp_output;
assign sign =a[n-1] ^ b[n-1];
localparam bias = 2**(m-1) -1;
assign expo_add= a[n-2:n-m-1] + b[n-2:n-m-1]; 
assign temp = expo_add - bias;
assign mant_mul = {1'b1,a[(n-m-2):0]} * {1'b1,b[(n-m-2):0]};
assign expo = mant_mul[2*(n-m)-1] ? temp+1:temp;
assign mant = mant_mul[2*(n-m)-1] ? mant_mul[(2*(n-m)-2):n-m] : mant_mul[(2*(n-m)-3):n-m-1];
assign temp_output={sign,expo[m-1:0],mant};

always@(*) 
    begin
    if(!a || !b ) begin
    out=0;
    overflow=0;
    underflow=0;
    end
   else if((~expo[m+1]&expo[m])||&expo[m-1:0]) begin
    overflow=1;
    underflow=0;
    out=0;
    end
   else if(expo[m+1]) begin
    underflow=1;
    overflow=0;
    out=0;
    end
   else begin
    out=temp_output;
    overflow=0;
    underflow=0;
    end
    
    end
endmodule
